module norgate(a,b,out);
input a,b;
output out;
nor a1(out,a,b);
endmodule