module notgate(a,out);
input a;
output out;
not a1(out,a);
endmodule